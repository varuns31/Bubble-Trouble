module fire_rom (
	input logic clock,
	input logic [9:0] address,
	output logic [8:0] q
);

logic [8:0] memory [0:543] /* synthesis ram_init_file = "./fire/fire.mif" */;

always_ff @ (posedge clock) begin
	q <= memory[address];
end

endmodule
