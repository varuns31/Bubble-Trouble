//module testbench();
//
//end
//endmodule
